*raw
    #include <parse.tab.h>

[a-z]+
    return IDENTIFIER;

*# vim: set sw=4 et:
