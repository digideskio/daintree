*raw
    #include <program.h>
    #include <parse.tab.h>
    #include <mem.h>

[a-z]+
    return IDENTIFIER;

*# vim: set sw=4 et:
